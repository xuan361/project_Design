module led(
    input CLK,
    input RESET,
    output [3:0] dig
    );




endmodule